library IEEE;
use IEEE.std_logic_1164.all;

--Entity
entity compressor is port
(
	X : in  std_logic;
	S : out std_logic
);
end entity;


-- Architecture
architecture logic of compressor is 
-- Signals


--Components

begin

end architecture;
