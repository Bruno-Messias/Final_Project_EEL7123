library IEEE;
use IEEE.std_logic_1164.all;

--Entity
entity compressor is port
(
	X : in  std_logic;
	S : out std_logic;
	s0: out std_logic_vector(3 downto 0)--teste 123
);
end entity;


-- Architecture
architecture logic of compressor is 
-- Signals


--Components

begin

end architecture;
